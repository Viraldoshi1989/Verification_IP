class config1;
	static mailbox #(txn) mbx=new();
endclass
